module ForwardingUnit (
    

    output  reg [1:0] FWD_rs1,
    output  reg [1:0] FWD_rs2
);
    
//------------------- parameter -------------------//    



endmodule
