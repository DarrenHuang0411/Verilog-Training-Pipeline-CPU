module ID_EXE_Reg (
    
    
    input   wire ID_pc;
    input   wire [32-1:0] rs1_data,
    input   wire [32-1:0] rs2_data,
    input   wire [6:0] funct7,
    input   wire [4:0] rs1_addr,
    input   wire [4:0] rs2_addr,
    input   wire [2:0] funct3,
    input   wire [4:0] rd_addr
);
    
endmodule
