module MEM_Stage (
    input   wire MEM_rd_sel,
    input   wire [:] MEM_DMread_sel,
    input   wire [:] MEM_DMwrite_sel,
);
    
    wire [:] MEM_rd_src;

endmodule
