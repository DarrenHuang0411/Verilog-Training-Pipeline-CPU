module Branch_Ctrl (
        
);
    
endmodule
