module IF_ID_Reg (

//Ctrl    
    input   wire HC_RW,
//I/O
    input   wire [32-1:0]   PC_in,
    input   wire [31:0]     instr_in,
    output  reg [32-1:0]    PC_ID_out,
    output  reg [31:0]      instr_out
);

reg [1:] ;

endmodule
