module ForwardingUnit (
    

    output  reg [:] FWDing2Mux2,
    output  reg [:] FWDing2Mux3

);
    
    



endmodule
