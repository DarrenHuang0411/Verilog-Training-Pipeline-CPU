`ifndef _PARAMETER_SETTING_
`define _PARAMETER_SETTING_

//DATA Parameter
    `define DATA_WIDTH      32

    `define OP_CODE         7
    `define FUNCTION_3      3
    `define FUNCTION_7      7

`endif