

module CLZ (
    input       [23:0]  significand_in,
    output  
);

    significand_s16
    significand_s16_8
    significand_s16_4
    significand_s16_2  
    
      
    m16
    m8
    m4
    m2
    m1
    always_comb begin
        if ((input && 0xff_ff00) == 0) begin
            
        end        
    end

endmodule